
//-----------------------------------Top_Processor_PMP ------------------------
// Top-level integration module for a single-cycle RISC-V processor
// augmented with Physical Memory Protection (PMP).
//
// This module serves as the system wrapper that:
//  - Connects the Control Unit and Datapath
//  - Routes decoded instruction fields to the controller
//  - Exposes internal signals for debugging and verification
//  - Aggregates PMP violations into meaningful system-level flags
//
// It represents the complete processor as observed by the testbench
// or verification environment.
//-------------------------------------------------------------------------------
`timescale 1ns / 1ps
`timescale 1ns / 1ps   // Duplicate timescale retained intentionally (no logic change)

module Top_Processor_PMP(
    input  wire        Clock,                     // System clock
    input  wire        Reset,                     // Global synchronous reset

    output wire [31:0] ALU_Result_Out,             // ALU result (debug/monitor)
    output wire [7:0]  PC_Out,                     // Current Program Counter
    output wire [6:0]  Opcode_Out,                 // Decoded instruction opcode
    output wire [2:0]  Funct3_Out,                 // Decoded funct3 field

    output wire        data_pmp_ok,                // Data access permission status
    output wire        instr_pmp_ok,               // Instruction fetch permission status

    // PMP violation visibility signals
    // These signals help distinguish the type of protection fault
    output wire        instr_exec_violation,       // Instruction execute violation
    output wire        data_read_violation,        // Data read violation
    output wire        data_write_violation,       // Data write violation
    output wire        PMP_Violation_Detected      // Aggregate PMP violation flag
);

    // ---------------- Control Signals ----------------
    // Generated by the Control Unit and consumed by the Datapath
    wire        Reg_Write;      // Register file write enable
    wire        ALU_Src;        // ALU operand source select
    wire [3:0]  ALU_CC;         // ALU control code
    wire        Mem_Read;       // Data memory read enable
    wire        Mem_Write;      // Data memory write enable
    wire        Mem_to_Reg;     // Write-back data select

    // ---------------- Instruction Fields ----------------
    // Extracted by the Datapath and fed back into the Control Unit
    wire [2:0]  Funct3;         // funct3 field
    wire [6:0]  Funct7;         // funct7 field
    wire [6:0]  Opcode;         // opcode field

    // ---------------- Datapath Result ----------------
    // ALU output exposed for debug and observation
    wire [31:0] Datapath_Result;

    // ---------------- Control Unit ----------------
    // Decodes instruction fields and generates high-level control signals
    Control_Unit control_unit (
        .opcode     (Opcode),
        .funct3     (Funct3),
        .funct7     (Funct7),
        .reg_write  (Reg_Write),
        .alu_src    (ALU_Src),
        .alu_cc     (ALU_CC),
        .mem_read   (Mem_Read),
        .mem_write  (Mem_Write),
        .mem_to_reg (Mem_to_Reg)
    );

    // ---------------- Datapath with PMP ----------------
    // Executes instructions, performs memory access,
    // and enforces PMP checks for both instruction fetch
    // and data memory access.
    Datapath_PMP datapath (
        .Clock           (Clock),
        .Reset           (Reset),
        .Reg_Write       (Reg_Write),
        .ALU_Src         (ALU_Src),
        .ALU_CC          (ALU_CC),
        .Mem_Read        (Mem_Read),
        .Mem_Write       (Mem_Write),
        .Mem_to_Reg      (Mem_to_Reg),
        .Funct3          (Funct3),
        .Funct7          (Funct7),
        .Opcode          (Opcode),
        .Datapath_Result (Datapath_Result),
        .data_pmp_ok     (data_pmp_ok),
        .instr_pmp_ok    (instr_pmp_ok),
        .PC              (PC_Out)
    );

    // ---------------- Output Assignments ----------------
    // Expose selected internal datapath signals
    assign ALU_Result_Out = Datapath_Result;
    assign Opcode_Out     = Opcode;
    assign Funct3_Out     = Funct3;

    // ---------------- PMP Violation Classification ----------------
    // These signals classify the type of PMP violation:
    // - Instruction execute violation: no execute permission
    // - Data read violation: load attempted without read permission
    // - Data write violation: store attempted without write permission
    assign instr_exec_violation = ~instr_pmp_ok;
    assign data_read_violation  = Mem_Read  & ~data_pmp_ok;
    assign data_write_violation = Mem_Write & ~data_pmp_ok;

    // ---------------- Global PMP Violation ----------------
    // Asserted whenever any type of PMP violation occurs.
    // Used as a system-level fault indication.
    assign PMP_Violation_Detected =
           instr_exec_violation |
           data_read_violation  |
           data_write_violation;

endmodule
